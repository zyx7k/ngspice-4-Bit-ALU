.subckt 3_OR nodeA nodeB nodeC output vdd gnd

X1 nodeA nodeB node1 vdd gnd OR
X2 nodeC node1 output vdd gnd OR

.ends 3_OR