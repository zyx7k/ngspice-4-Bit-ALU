.subckt AND_BLOCK A0 A1 A2 A3 B0 B1 B2 B3 AB_0 AB_1 AB_2 AB_3 vdd gnd

X1 A0 B0 AB_0 vdd gnd AND
X2 A1 B1 AB_1 vdd gnd AND
X3 A2 B2 AB_2 vdd gnd AND
X4 A3 B3 AB_3 vdd gnd AND

.ends AND_BLOCK