.subckt 5_AND nodeA nodeB nodeC nodeD nodeE output vdd gnd

X1 nodeA nodeB nodeC nodeD node1 vdd gnd 4_AND
X2 nodeE node1 output vdd gnd AND

.ends 5_AND