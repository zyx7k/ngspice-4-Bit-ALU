.subckt ENABLE E A0 A1 A2 A3 B0 B1 B2 B3 A0_E A1_E A2_E A3_E B0_E B1_E B2_E B3_E vdd gnd 

X1 A0 E A0_E vdd gnd AND
X2 A1 E A1_E vdd gnd AND
X3 A2 E A2_E vdd gnd AND
X4 A3 E A3_E vdd gnd AND

X5 B0 E B0_E vdd gnd AND
X6 B1 E B1_E vdd gnd AND
X7 B2 E B2_E vdd gnd AND
X8 B3 E B3_E vdd gnd AND

.ends ENABLE    