.subckt 4_AND nodeA nodeB nodeC nodeD output vdd gnd

X1 nodeA nodeB nodeC node1 vdd gnd 3_AND
X2 nodeD node1 output vdd gnd AND

.ends 4_AND