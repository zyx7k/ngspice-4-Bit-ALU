.subckt 4_OR nodeA nodeB nodeC nodeD output vdd gnd

X1 nodeA nodeB nodeC node1 vdd gnd 3_OR
X2 nodeD node1 output vdd gnd OR

.ends 4_OR